`timescale 1ns / 1ps

module jit_switch #(
  parameter integer NUM_ACCs = 2
)
(
  output  wire             sCMD_tready ,
  input   wire             sCMD_tvalid ,
  input   wire  [31 : 0]   sCMD_tdata  ,

//input   wire             mRSP_tready ,
//output  wire             mRSP_tvalid ,
//output  wire  [31 : 0]   mRSP_tdata  ,
//// -----------------------------------
  output  wire             s1A_tready  ,
  input   wire             s1A_tvalid  ,
  input   wire  [31 : 0]   s1A_tdata   ,

  output  wire             s1B_tready  ,
  input   wire             s1B_tvalid  ,
  input   wire  [31 : 0]   s1B_tdata   ,

  input   wire             m1C_tready  ,
  output  wire             m1C_tvalid  ,
  output  wire  [31 : 0]   m1C_tdata   ,

  output  wire             s1AT_tready ,
  input   wire             s1AT_tvalid ,
  input   wire  [31 : 0]   s1AT_tdata  ,

  output  wire             s1BT_tready ,
  input   wire             s1BT_tvalid ,
  input   wire  [31 : 0]   s1BT_tdata  ,

  input   wire             m1CT_tready ,
  output  wire             m1CT_tvalid ,
  output  wire  [31 : 0]   m1CT_tdata  ,

  output  wire             s1C_tready  ,
  input   wire             s1C_tvalid  ,
  input   wire  [31 : 0]   s1C_tdata   ,

  input   wire             m1A_tready  ,
  output  wire             m1A_tvalid  ,
  output  wire  [31 : 0]   m1A_tdata   ,

  input   wire             m1B_tready  ,
  output  wire             m1B_tvalid  ,
  output  wire  [31 : 0]   m1B_tdata   ,
  // -----------------------------------
  output  wire             s2A_tready  ,
  input   wire             s2A_tvalid  ,
  input   wire  [31 : 0]   s2A_tdata   ,

  output  wire             s2B_tready  ,
  input   wire             s2B_tvalid  ,
  input   wire  [31 : 0]   s2B_tdata   ,

  input   wire             m2C_tready  ,
  output  wire             m2C_tvalid  ,
  output  wire  [31 : 0]   m2C_tdata   ,

  output  wire             s2AT_tready ,
  input   wire             s2AT_tvalid ,
  input   wire  [31 : 0]   s2AT_tdata  ,

  output  wire             s2BT_tready ,
  input   wire             s2BT_tvalid ,
  input   wire  [31 : 0]   s2BT_tdata  ,

  input   wire             m2CT_tready ,
  output  wire             m2CT_tvalid ,
  output  wire  [31 : 0]   m2CT_tdata  ,

  output  wire             s2C_tready  ,
  input   wire             s2C_tvalid  ,
  input   wire  [31 : 0]   s2C_tdata   ,

  input   wire             m2A_tready  ,
  output  wire             m2A_tvalid  ,
  output  wire  [31 : 0]   m2A_tdata   ,

  input   wire             m2B_tready  ,
  output  wire             m2B_tvalid  ,
  output  wire  [31 : 0]   m2B_tdata   ,
  // -----------------------------------
  output  wire             s3A_tready  ,
  input   wire             s3A_tvalid  ,
  input   wire  [31 : 0]   s3A_tdata   ,

  output  wire             s3B_tready  ,
  input   wire             s3B_tvalid  ,
  input   wire  [31 : 0]   s3B_tdata   ,

  input   wire             m3C_tready  ,
  output  wire             m3C_tvalid  ,
  output  wire  [31 : 0]   m3C_tdata   ,

  output  wire             s3AT_tready ,
  input   wire             s3AT_tvalid ,
  input   wire  [31 : 0]   s3AT_tdata  ,

  output  wire             s3BT_tready ,
  input   wire             s3BT_tvalid ,
  input   wire  [31 : 0]   s3BT_tdata  ,

  input   wire             m3CT_tready ,
  output  wire             m3CT_tvalid ,
  output  wire  [31 : 0]   m3CT_tdata  ,

  output  wire             s3C_tready  ,
  input   wire             s3C_tvalid  ,
  input   wire  [31 : 0]   s3C_tdata   ,

  input   wire             m3A_tready  ,
  output  wire             m3A_tvalid  ,
  output  wire  [31 : 0]   m3A_tdata   ,

  input   wire             m3B_tready  ,
  output  wire             m3B_tvalid  ,
  output  wire  [31 : 0]   m3B_tdata   ,
  // -----------------------------------
  output  wire             s4A_tready  ,
  input   wire             s4A_tvalid  ,
  input   wire  [31 : 0]   s4A_tdata   ,

  output  wire             s4B_tready  ,
  input   wire             s4B_tvalid  ,
  input   wire  [31 : 0]   s4B_tdata   ,

  input   wire             m4C_tready  ,
  output  wire             m4C_tvalid  ,
  output  wire  [31 : 0]   m4C_tdata   ,

  output  wire             s4AT_tready ,
  input   wire             s4AT_tvalid ,
  input   wire  [31 : 0]   s4AT_tdata  ,

  output  wire             s4BT_tready ,
  input   wire             s4BT_tvalid ,
  input   wire  [31 : 0]   s4BT_tdata  ,

  input   wire             m4CT_tready ,
  output  wire             m4CT_tvalid ,
  output  wire  [31 : 0]   m4CT_tdata  ,

  output  wire             s4C_tready  ,
  input   wire             s4C_tvalid  ,
  input   wire  [31 : 0]   s4C_tdata   ,

  input   wire             m4A_tready  ,
  output  wire             m4A_tvalid  ,
  output  wire  [31 : 0]   m4A_tdata   ,

  input   wire             m4B_tready  ,
  output  wire             m4B_tvalid  ,
  output  wire  [31 : 0]   m4B_tdata   ,
  // -----------------------------------
  output  wire             s5A_tready  ,
  input   wire             s5A_tvalid  ,
  input   wire  [31 : 0]   s5A_tdata   ,

  output  wire             s5B_tready  ,
  input   wire             s5B_tvalid  ,
  input   wire  [31 : 0]   s5B_tdata   ,

  input   wire             m5C_tready  ,
  output  wire             m5C_tvalid  ,
  output  wire  [31 : 0]   m5C_tdata   ,

  output  wire             s5AT_tready ,
  input   wire             s5AT_tvalid ,
  input   wire  [31 : 0]   s5AT_tdata  ,

  output  wire             s5BT_tready ,
  input   wire             s5BT_tvalid ,
  input   wire  [31 : 0]   s5BT_tdata  ,

  input   wire             m5CT_tready ,
  output  wire             m5CT_tvalid ,
  output  wire  [31 : 0]   m5CT_tdata  ,

  output  wire             s5C_tready  ,
  input   wire             s5C_tvalid  ,
  input   wire  [31 : 0]   s5C_tdata   ,

  input   wire             m5A_tready  ,
  output  wire             m5A_tvalid  ,
  output  wire  [31 : 0]   m5A_tdata   ,

  input   wire             m5B_tready  ,
  output  wire             m5B_tvalid  ,
  output  wire  [31 : 0]   m5B_tdata   ,
  // -----------------------------------
  output  wire             s6A_tready  ,
  input   wire             s6A_tvalid  ,
  input   wire  [31 : 0]   s6A_tdata   ,

  output  wire             s6B_tready  ,
  input   wire             s6B_tvalid  ,
  input   wire  [31 : 0]   s6B_tdata   ,

  input   wire             m6C_tready  ,
  output  wire             m6C_tvalid  ,
  output  wire  [31 : 0]   m6C_tdata   ,

  output  wire             s6AT_tready ,
  input   wire             s6AT_tvalid ,
  input   wire  [31 : 0]   s6AT_tdata  ,

  output  wire             s6BT_tready ,
  input   wire             s6BT_tvalid ,
  input   wire  [31 : 0]   s6BT_tdata  ,

  input   wire             m6CT_tready ,
  output  wire             m6CT_tvalid ,
  output  wire  [31 : 0]   m6CT_tdata  ,

  output  wire             s6C_tready  ,
  input   wire             s6C_tvalid  ,
  input   wire  [31 : 0]   s6C_tdata   ,

  input   wire             m6A_tready  ,
  output  wire             m6A_tvalid  ,
  output  wire  [31 : 0]   m6A_tdata   ,

  input   wire             m6B_tready  ,
  output  wire             m6B_tvalid  ,
  output  wire  [31 : 0]   m6B_tdata   ,
  // -----------------------------------
  output  wire             s7A_tready  ,
  input   wire             s7A_tvalid  ,
  input   wire  [31 : 0]   s7A_tdata   ,

  output  wire             s7B_tready  ,
  input   wire             s7B_tvalid  ,
  input   wire  [31 : 0]   s7B_tdata   ,

  input   wire             m7C_tready  ,
  output  wire             m7C_tvalid  ,
  output  wire  [31 : 0]   m7C_tdata   ,

  output  wire             s7AT_tready ,
  input   wire             s7AT_tvalid ,
  input   wire  [31 : 0]   s7AT_tdata  ,

  output  wire             s7BT_tready ,
  input   wire             s7BT_tvalid ,
  input   wire  [31 : 0]   s7BT_tdata  ,

  input   wire             m7CT_tready ,
  output  wire             m7CT_tvalid ,
  output  wire  [31 : 0]   m7CT_tdata  ,

  output  wire             s7C_tready  ,
  input   wire             s7C_tvalid  ,
  input   wire  [31 : 0]   s7C_tdata   ,

  input   wire             m7A_tready  ,
  output  wire             m7A_tvalid  ,
  output  wire  [31 : 0]   m7A_tdata   ,

  input   wire             m7B_tready  ,
  output  wire             m7B_tvalid  ,
  output  wire  [31 : 0]   m7B_tdata   ,
  // -----------------------------------
  output  wire             s8A_tready  ,
  input   wire             s8A_tvalid  ,
  input   wire  [31 : 0]   s8A_tdata   ,

  output  wire             s8B_tready  ,
  input   wire             s8B_tvalid  ,
  input   wire  [31 : 0]   s8B_tdata   ,

  input   wire             m8C_tready  ,
  output  wire             m8C_tvalid  ,
  output  wire  [31 : 0]   m8C_tdata   ,

  output  wire             s8AT_tready ,
  input   wire             s8AT_tvalid ,
  input   wire  [31 : 0]   s8AT_tdata  ,

  output  wire             s8BT_tready ,
  input   wire             s8BT_tvalid ,
  input   wire  [31 : 0]   s8BT_tdata  ,

  input   wire             m8CT_tready ,
  output  wire             m8CT_tvalid ,
  output  wire  [31 : 0]   m8CT_tdata  ,

  output  wire             s8C_tready  ,
  input   wire             s8C_tvalid  ,
  input   wire  [31 : 0]   s8C_tdata   ,

  input   wire             m8A_tready  ,
  output  wire             m8A_tvalid  ,
  output  wire  [31 : 0]   m8A_tdata   ,

  input   wire             m8B_tready  ,
  output  wire             m8B_tvalid  ,
  output  wire  [31 : 0]   m8B_tdata   ,
//// -----------------------------------
//input   wire             ap1_done    ,
//input   wire             ap1_idle    ,
//input   wire             ap1_ready   ,
//output  wire             ap1_start   ,
  output  wire  [15 : 0]   ap1_arg1_V  ,
  output  wire  [15 : 0]   ap1_arg2_V  ,
  output  wire  [15 : 0]   ap1_arg3_V  ,
//// -----------------------------------
//input   wire             ap2_done    ,
//input   wire             ap2_idle    ,
//input   wire             ap2_ready   ,
//output  wire             ap2_start   ,
  output  wire  [15 : 0]   ap2_arg1_V  ,
  output  wire  [15 : 0]   ap2_arg2_V  ,
  output  wire  [15 : 0]   ap2_arg3_V  ,
//// -----------------------------------
//input   wire             ap3_done    ,
//input   wire             ap3_idle    ,
//input   wire             ap3_ready   ,
//output  wire             ap3_start   ,
  output  wire  [15 : 0]   ap3_arg1_V  ,
  output  wire  [15 : 0]   ap3_arg2_V  ,
  output  wire  [15 : 0]   ap3_arg3_V  ,
//// -----------------------------------
//input   wire             ap4_done    ,
//input   wire             ap4_idle    ,
//input   wire             ap4_ready   ,
//output  wire             ap4_start   ,
  output  wire  [15 : 0]   ap4_arg1_V  ,
  output  wire  [15 : 0]   ap4_arg2_V  ,
  output  wire  [15 : 0]   ap4_arg3_V  ,
//// -----------------------------------
//input   wire             ap5_done    ,
//input   wire             ap5_idle    ,
//input   wire             ap5_ready   ,
//output  wire             ap5_start   ,
  output  wire  [15 : 0]   ap5_arg1_V  ,
  output  wire  [15 : 0]   ap5_arg2_V  ,
  output  wire  [15 : 0]   ap5_arg3_V  ,
//// -----------------------------------
//input   wire             ap6_done    ,
//input   wire             ap6_idle    ,
//input   wire             ap6_ready   ,
//output  wire             ap6_start   ,
  output  wire  [15 : 0]   ap6_arg1_V  ,
  output  wire  [15 : 0]   ap6_arg2_V  ,
  output  wire  [15 : 0]   ap6_arg3_V  ,
//// -----------------------------------
//input   wire             ap7_done    ,
//input   wire             ap7_idle    ,
//input   wire             ap7_ready   ,
//output  wire             ap7_start   ,
  output  wire  [15 : 0]   ap7_arg1_V  ,
  output  wire  [15 : 0]   ap7_arg2_V  ,
  output  wire  [15 : 0]   ap7_arg3_V  ,
//// -----------------------------------
//input   wire             ap8_done    ,
//input   wire             ap8_idle    ,
//input   wire             ap8_ready   ,
//output  wire             ap8_start   ,
  output  wire  [15 : 0]   ap8_arg1_V  ,
  output  wire  [15 : 0]   ap8_arg2_V  ,
  output  wire  [15 : 0]   ap8_arg3_V  ,
  // -----------------------------------
  input   wire             ACLK        ,
  input   wire             ARESETN
);
  wire             w1cA_tready  ;
  wire             w1cA_tvalid  ;
  wire  [31 : 0]   w1cA_tdata   ;
  wire             w1cB_tready  ;
  wire             w1cB_tvalid  ;
  wire  [31 : 0]   w1cB_tdata   ;
  wire             w1cC_tready  ;
  wire             w1cC_tvalid  ;
  wire  [31 : 0]   w1cC_tdata   ;

  wire             w2cA_tready  ;
  wire             w2cA_tvalid  ;
  wire  [31 : 0]   w2cA_tdata   ;
  wire             w2cB_tready  ;
  wire             w2cB_tvalid  ;
  wire  [31 : 0]   w2cB_tdata   ;
  wire             w2cC_tready  ;
  wire             w2cC_tvalid  ;
  wire  [31 : 0]   w2cC_tdata   ;

  wire             w3cA_tready  ;
  wire             w3cA_tvalid  ;
  wire  [31 : 0]   w3cA_tdata   ;
  wire             w3cB_tready  ;
  wire             w3cB_tvalid  ;
  wire  [31 : 0]   w3cB_tdata   ;
  wire             w3cC_tready  ;
  wire             w3cC_tvalid  ;
  wire  [31 : 0]   w3cC_tdata   ;

  wire             w4cA_tready  ;
  wire             w4cA_tvalid  ;
  wire  [31 : 0]   w4cA_tdata   ;
  wire             w4cB_tready  ;
  wire             w4cB_tvalid  ;
  wire  [31 : 0]   w4cB_tdata   ;
  wire             w4cC_tready  ;
  wire             w4cC_tvalid  ;
  wire  [31 : 0]   w4cC_tdata   ;

  wire             w5cA_tready  ;
  wire             w5cA_tvalid  ;
  wire  [31 : 0]   w5cA_tdata   ;
  wire             w5cB_tready  ;
  wire             w5cB_tvalid  ;
  wire  [31 : 0]   w5cB_tdata   ;
  wire             w5cC_tready  ;
  wire             w5cC_tvalid  ;
  wire  [31 : 0]   w5cC_tdata   ;

  wire             w6cA_tready  ;
  wire             w6cA_tvalid  ;
  wire  [31 : 0]   w6cA_tdata   ;
  wire             w6cB_tready  ;
  wire             w6cB_tvalid  ;
  wire  [31 : 0]   w6cB_tdata   ;
  wire             w6cC_tready  ;
  wire             w6cC_tvalid  ;
  wire  [31 : 0]   w6cC_tdata   ;

  wire             w7cA_tready  ;
  wire             w7cA_tvalid  ;
  wire  [31 : 0]   w7cA_tdata   ;
  wire             w7cB_tready  ;
  wire             w7cB_tvalid  ;
  wire  [31 : 0]   w7cB_tdata   ;
  wire             w7cC_tready  ;
  wire             w7cC_tvalid  ;
  wire  [31 : 0]   w7cC_tdata   ;

  wire             w8cA_tready  ;
  wire             w8cA_tvalid  ;
  wire  [31 : 0]   w8cA_tdata   ;
  wire             w8cB_tready  ;
  wire             w8cB_tvalid  ;
  wire  [31 : 0]   w8cB_tdata   ;
  wire             w8cC_tready  ;
  wire             w8cC_tvalid  ;
  wire  [31 : 0]   w8cC_tdata   ;

  wire  [ 3 : 0]   acc1_A1      ;
  wire  [ 3 : 0]   acc1_B1      ;
  wire  [ 5 : 0]   acc1_C1      ;
  wire  [ 3 : 0]   acc2_A1      ;
  wire  [ 3 : 0]   acc2_B1      ;
  wire  [ 5 : 0]   acc2_C1      ;
  wire  [ 3 : 0]   acc3_A1      ;
  wire  [ 3 : 0]   acc3_B1      ;
  wire  [ 5 : 0]   acc3_C1      ;
  wire  [ 3 : 0]   acc4_A1      ;
  wire  [ 3 : 0]   acc4_B1      ;
  wire  [ 5 : 0]   acc4_C1      ;
  wire  [ 3 : 0]   acc5_A1      ;
  wire  [ 3 : 0]   acc5_B1      ;
  wire  [ 5 : 0]   acc5_C1      ;
  wire  [ 3 : 0]   acc6_A1      ;
  wire  [ 3 : 0]   acc6_B1      ;
  wire  [ 5 : 0]   acc6_C1      ;
  wire  [ 3 : 0]   acc7_A1      ;
  wire  [ 3 : 0]   acc7_B1      ;
  wire  [ 5 : 0]   acc7_C1      ;
  wire  [ 3 : 0]   acc8_A1      ;
  wire  [ 3 : 0]   acc8_B1      ;
  wire  [ 5 : 0]   acc8_C1      ;
//       _    ____ ____           ____
//      / \  / ___/ ___|___   _  |___ \
//     / _ \| |  | |   / __| (_)   __) |
//    / ___ \ |__| |___\__ \  _   / __/
//   /_/   \_\____\____|___/ (_) |_____|
//
generate if (NUM_ACCs == 2) begin

  jit_couple u_acc1_couple (
    .sInA_tready      (s1A_tready   ),
    .sInA_tvalid      (s1A_tvalid   ),
    .sInA_tdata       (s1A_tdata    ),
    .sInB_tready      (s1B_tready   ),
    .sInB_tvalid      (s1B_tvalid   ),
    .sInB_tdata       (s1B_tdata    ),
    .mOutC_tready     (m1C_tready   ),
    .mOutC_tvalid     (m1C_tvalid   ),
    .mOutC_tdata      (m1C_tdata    ),
    .sInAT_tready     (s1AT_tready  ),
    .sInAT_tvalid     (s1AT_tvalid  ),
    .sInAT_tdata      (s1AT_tdata   ),
    .sInBT_tready     (s1BT_tready  ),
    .sInBT_tvalid     (s1BT_tvalid  ),
    .sInBT_tdata      (s1BT_tdata   ),
    .mOutCT_tready    (m1CT_tready  ),
    .mOutCT_tvalid    (m1CT_tvalid  ),
    .mOutCT_tdata     (m1CT_tdata   ),
    .scInA_tready     (w1cA_tready  ),
    .scInA_tvalid     (w1cA_tvalid  ),
    .scInA_tdata      (w1cA_tdata   ),
    .scInB_tready     (w1cB_tready  ),
    .scInB_tvalid     (w1cB_tvalid  ),
    .scInB_tdata      (w1cB_tdata   ),
    .mcOutC_tready    (w1cC_tready  ),
    .mcOutC_tvalid    (w1cC_tvalid  ),
    .mcOutC_tdata     (w1cC_tdata   ),
    .sAccInC_tready   (s1C_tready   ),
    .sAccInC_tvalid   (s1C_tvalid   ),
    .sAccInC_tdata    (s1C_tdata    ),
    .mAccOutA_tready  (m1A_tready   ),
    .mAccOutA_tvalid  (m1A_tvalid   ),
    .mAccOutA_tdata   (m1A_tdata    ),
    .mAccOutB_tready  (m1B_tready   ),
    .mAccOutB_tvalid  (m1B_tvalid   ),
    .mAccOutB_tdata   (m1B_tdata    ),
    .CONF             (acc1_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc2_couple (
    .sInA_tready      (s2A_tready   ),
    .sInA_tvalid      (s2A_tvalid   ),
    .sInA_tdata       (s2A_tdata    ),
    .sInB_tready      (s2B_tready   ),
    .sInB_tvalid      (s2B_tvalid   ),
    .sInB_tdata       (s2B_tdata    ),
    .mOutC_tready     (m2C_tready   ),
    .mOutC_tvalid     (m2C_tvalid   ),
    .mOutC_tdata      (m2C_tdata    ),
    .sInAT_tready     (s2AT_tready  ),
    .sInAT_tvalid     (s2AT_tvalid  ),
    .sInAT_tdata      (s2AT_tdata   ),
    .sInBT_tready     (s2BT_tready  ),
    .sInBT_tvalid     (s2BT_tvalid  ),
    .sInBT_tdata      (s2BT_tdata   ),
    .mOutCT_tready    (m2CT_tready  ),
    .mOutCT_tvalid    (m2CT_tvalid  ),
    .mOutCT_tdata     (m2CT_tdata   ),
    .scInA_tready     (w2cA_tready  ),
    .scInA_tvalid     (w2cA_tvalid  ),
    .scInA_tdata      (w2cA_tdata   ),
    .scInB_tready     (w2cB_tready  ),
    .scInB_tvalid     (w2cB_tvalid  ),
    .scInB_tdata      (w2cB_tdata   ),
    .mcOutC_tready    (w2cC_tready  ),
    .mcOutC_tvalid    (w2cC_tvalid  ),
    .mcOutC_tdata     (w2cC_tdata   ),
    .sAccInC_tready   (s2C_tready   ),
    .sAccInC_tvalid   (s2C_tvalid   ),
    .sAccInC_tdata    (s2C_tdata    ),
    .mAccOutA_tready  (m2A_tready   ),
    .mAccOutA_tvalid  (m2A_tvalid   ),
    .mAccOutA_tdata   (m2A_tdata    ),
    .mAccOutB_tready  (m2B_tready   ),
    .mAccOutB_tvalid  (m2B_tvalid   ),
    .mAccOutB_tdata   (m2B_tdata    ),
    .CONF             (acc2_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_crossbar #(NUM_ACCs) u_crossbar (
    .CONF1_A       (acc1_A1         ),
    .CONF1_B       (acc1_B1         ),
    .sC1_tready    (w1cC_tready     ),
    .sC1_tvalid    (w1cC_tvalid     ),
    .sC1_tdata     (w1cC_tdata      ),
    .mA1_tready    (w1cA_tready     ),
    .mA1_tvalid    (w1cA_tvalid     ),
    .mA1_tdata     (w1cA_tdata      ),
    .mB1_tready    (w1cB_tready     ),
    .mB1_tvalid    (w1cB_tvalid     ),
    .mB1_tdata     (w1cB_tdata      ),
    .CONF2_A       (acc2_A1         ),
    .CONF2_B       (acc2_B1         ),
    .sC2_tready    (w2cC_tready     ),
    .sC2_tvalid    (w2cC_tvalid     ),
    .sC2_tdata     (w2cC_tdata      ),
    .mA2_tready    (w2cA_tready     ),
    .mA2_tvalid    (w2cA_tvalid     ),
    .mA2_tdata     (w2cA_tdata      ),
    .mB2_tready    (w2cB_tready     ),
    .mB2_tvalid    (w2cB_tvalid     ),
    .mB2_tdata     (w2cB_tdata      ),
    .CONF3_A       (acc3_A1         ),
    .CONF3_B       (acc3_B1         ),
    .sC3_tready    (w3cC_tready     ),
    .sC3_tvalid    ( 1'd0           ),
    .sC3_tdata     (32'd0           ),
    .mA3_tready    ( 1'd0           ),
    .mA3_tvalid    (w3cA_tvalid     ),
    .mA3_tdata     (w3cA_tdata      ),
    .mB3_tready    ( 1'd0           ),
    .mB3_tvalid    (w3cB_tvalid     ),
    .mB3_tdata     (w3cB_tdata      ),
    .CONF4_A       (acc4_A1         ),
    .CONF4_B       (acc4_B1         ),
    .sC4_tready    (w4cC_tready     ),
    .sC4_tvalid    ( 1'd0           ),
    .sC4_tdata     (32'd0           ),
    .mA4_tready    ( 1'd0           ),
    .mA4_tvalid    (w4cA_tvalid     ),
    .mA4_tdata     (w4cA_tdata      ),
    .mB4_tready    ( 1'd0           ),
    .mB4_tvalid    (w4cB_tvalid     ),
    .mB4_tdata     (w4cB_tdata      ),
    .CONF5_A       (acc5_A1         ),
    .CONF5_B       (acc5_B1         ),
    .sC5_tready    (w5cC_tready     ),
    .sC5_tvalid    ( 1'd0           ),
    .sC5_tdata     (32'd0           ),
    .mA5_tready    ( 1'd0           ),
    .mA5_tvalid    (w5cA_tvalid     ),
    .mA5_tdata     (w5cA_tdata      ),
    .mB5_tready    ( 1'd0           ),
    .mB5_tvalid    (w5cB_tvalid     ),
    .mB5_tdata     (w5cB_tdata      ),
    .CONF6_A       (acc6_A1         ),
    .CONF6_B       (acc6_B1         ),
    .sC6_tready    (w6cC_tready     ),
    .sC6_tvalid    ( 1'd0           ),
    .sC6_tdata     (32'd0           ),
    .mA6_tready    ( 1'd0           ),
    .mA6_tvalid    (w6cA_tvalid     ),
    .mA6_tdata     (w6cA_tdata      ),
    .mB6_tready    ( 1'd0           ),
    .mB6_tvalid    (w6cB_tvalid     ),
    .mB6_tdata     (w6cB_tdata      ),
    .CONF7_A       (acc7_A1         ),
    .CONF7_B       (acc7_B1         ),
    .sC7_tready    (w7cC_tready     ),
    .sC7_tvalid    ( 1'd0           ),
    .sC7_tdata     (32'd0           ),
    .mA7_tready    ( 1'd0           ),
    .mA7_tvalid    (w7cA_tvalid     ),
    .mA7_tdata     (w7cA_tdata      ),
    .mB7_tready    ( 1'd0           ),
    .mB7_tvalid    (w7cB_tvalid     ),
    .mB7_tdata     (w7cB_tdata      ),
    .CONF8_A       (acc8_A1         ),
    .CONF8_B       (acc8_B1         ),
    .sC8_tready    (w8cC_tready     ),
    .sC8_tvalid    ( 1'd0           ),
    .sC8_tdata     (32'd0           ),
    .mA8_tready    ( 1'd0           ),
    .mA8_tvalid    (w8cA_tvalid     ),
    .mA8_tdata     (w8cA_tdata      ),
    .mB8_tready    ( 1'd0           ),
    .mB8_tvalid    (w8cB_tvalid     ),
    .mB8_tdata     (w8cB_tdata      ),
    .ACLK          (ACLK            ),
    .ARESETN       (ARESETN         )
  );

  jit_dispatch #(NUM_ACCs) u_dispatch(
    .sR_tready     (sCMD_tready     ),
    .sR_tvalid     (sCMD_tvalid     ),
    .sR_tdata      (sCMD_tdata      ),
//  .mR_tready     (mRSP_tready     ),
//  .mR_tvalid     (mRSP_tvalid     ),
//  .mR_tdata      (mRSP_tdata      ),
    .acc1_A1       (acc1_A1         ),
    .acc1_B1       (acc1_B1         ),
    .acc1_C1       (acc1_C1         ),
    .acc1_R1       (ap1_arg1_V      ),
    .acc1_R2       (ap1_arg2_V      ),
    .acc1_R3       (ap1_arg3_V      ),
//  .acc1_done     (ap1_done        ),
//  .acc1_idle     (ap1_idle        ),
//  .acc1_ready    (ap1_ready       ),
//  .acc1_start    (ap1_start       ),
    .acc2_A1       (acc2_A1         ),
    .acc2_B1       (acc2_B1         ),
    .acc2_C1       (acc2_C1         ),
    .acc2_R1       (ap2_arg1_V      ),
    .acc2_R2       (ap2_arg2_V      ),
    .acc2_R3       (ap2_arg3_V      ),
//  .acc2_done     (ap2_done        ),
//  .acc2_idle     (ap2_idle        ),
//  .acc2_ready    (ap2_ready       ),
//  .acc2_start    (ap2_start       ),
    .acc3_A1       (acc3_A1         ),
    .acc3_B1       (acc3_B1         ),
    .acc3_C1       (acc3_C1         ),
    .acc3_R1       (ap3_arg1_V      ),
    .acc3_R2       (ap3_arg2_V      ),
    .acc3_R3       (ap3_arg3_V      ),
//  .acc3_done     (ap3_done        ),
//  .acc3_idle     (ap3_idle        ),
//  .acc3_ready    (ap3_ready       ),
//  .acc3_start    (ap3_start       ),
    .acc4_A1       (acc4_A1         ),
    .acc4_B1       (acc4_B1         ),
    .acc4_C1       (acc4_C1         ),
    .acc4_R1       (ap4_arg1_V      ),
    .acc4_R2       (ap4_arg2_V      ),
    .acc4_R3       (ap4_arg3_V      ),
//  .acc4_done     (ap4_done        ),
//  .acc4_idle     (ap4_idle        ),
//  .acc4_ready    (ap4_ready       ),
//  .acc4_start    (ap4_start       ),
    .acc5_A1       (acc5_A1         ),
    .acc5_B1       (acc5_B1         ),
    .acc5_C1       (acc5_C1         ),
    .acc5_R1       (ap5_arg1_V      ),
    .acc5_R2       (ap5_arg2_V      ),
    .acc5_R3       (ap5_arg3_V      ),
//  .acc5_done     (ap5_done        ),
//  .acc5_idle     (ap5_idle        ),
//  .acc5_ready    (ap5_ready       ),
//  .acc5_start    (ap5_start       ),
    .acc6_A1       (acc6_A1         ),
    .acc6_B1       (acc6_B1         ),
    .acc6_C1       (acc6_C1         ),
    .acc6_R1       (ap6_arg1_V      ),
    .acc6_R2       (ap6_arg2_V      ),
    .acc6_R3       (ap6_arg3_V      ),
//  .acc6_done     (ap6_done        ),
//  .acc6_idle     (ap6_idle        ),
//  .acc6_ready    (ap6_ready       ),
//  .acc6_start    (ap6_start       ),
    .acc7_A1       (acc7_A1         ),
    .acc7_B1       (acc7_B1         ),
    .acc7_C1       (acc7_C1         ),
    .acc7_R1       (ap7_arg1_V      ),
    .acc7_R2       (ap7_arg2_V      ),
    .acc7_R3       (ap7_arg3_V      ),
//  .acc7_done     (ap7_done        ),
//  .acc7_idle     (ap7_idle        ),
//  .acc7_ready    (ap7_ready       ),
//  .acc7_start    (ap7_start       ),
    .acc8_A1       (acc8_A1         ),
    .acc8_B1       (acc8_B1         ),
    .acc8_C1       (acc8_C1         ),
    .acc8_R1       (ap8_arg1_V      ),
    .acc8_R2       (ap8_arg2_V      ),
    .acc8_R3       (ap8_arg3_V      ),
//  .acc8_done     (ap8_done        ),
//  .acc8_idle     (ap8_idle        ),
//  .acc8_ready    (ap8_ready       ),
//  .acc8_start    (ap8_start       ),
    .ACLK          (ACLK            ),
    .ARESETN       (ARESETN         )
  );

end
endgenerate // NUM_ACCs == 2

//       _    ____ ____           _  _
//      / \  / ___/ ___|___   _  | || |
//     / _ \| |  | |   / __| (_) | || |_
//    / ___ \ |__| |___\__ \  _  |__   _|
//   /_/   \_\____\____|___/ (_)    |_|
//
generate if (NUM_ACCs == 4) begin

  jit_couple u_acc1_couple (
    .sInA_tready      (s1A_tready   ),
    .sInA_tvalid      (s1A_tvalid   ),
    .sInA_tdata       (s1A_tdata    ),
    .sInB_tready      (s1B_tready   ),
    .sInB_tvalid      (s1B_tvalid   ),
    .sInB_tdata       (s1B_tdata    ),
    .mOutC_tready     (m1C_tready   ),
    .mOutC_tvalid     (m1C_tvalid   ),
    .mOutC_tdata      (m1C_tdata    ),
    .sInAT_tready     (s1AT_tready  ),
    .sInAT_tvalid     (s1AT_tvalid  ),
    .sInAT_tdata      (s1AT_tdata   ),
    .sInBT_tready     (s1BT_tready  ),
    .sInBT_tvalid     (s1BT_tvalid  ),
    .sInBT_tdata      (s1BT_tdata   ),
    .mOutCT_tready    (m1CT_tready  ),
    .mOutCT_tvalid    (m1CT_tvalid  ),
    .mOutCT_tdata     (m1CT_tdata   ),
    .scInA_tready     (w1cA_tready  ),
    .scInA_tvalid     (w1cA_tvalid  ),
    .scInA_tdata      (w1cA_tdata   ),
    .scInB_tready     (w1cB_tready  ),
    .scInB_tvalid     (w1cB_tvalid  ),
    .scInB_tdata      (w1cB_tdata   ),
    .mcOutC_tready    (w1cC_tready  ),
    .mcOutC_tvalid    (w1cC_tvalid  ),
    .mcOutC_tdata     (w1cC_tdata   ),
    .sAccInC_tready   (s1C_tready   ),
    .sAccInC_tvalid   (s1C_tvalid   ),
    .sAccInC_tdata    (s1C_tdata    ),
    .mAccOutA_tready  (m1A_tready   ),
    .mAccOutA_tvalid  (m1A_tvalid   ),
    .mAccOutA_tdata   (m1A_tdata    ),
    .mAccOutB_tready  (m1B_tready   ),
    .mAccOutB_tvalid  (m1B_tvalid   ),
    .mAccOutB_tdata   (m1B_tdata    ),
    .CONF             (acc1_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc2_couple (
    .sInA_tready      (s2A_tready   ),
    .sInA_tvalid      (s2A_tvalid   ),
    .sInA_tdata       (s2A_tdata    ),
    .sInB_tready      (s2B_tready   ),
    .sInB_tvalid      (s2B_tvalid   ),
    .sInB_tdata       (s2B_tdata    ),
    .mOutC_tready     (m2C_tready   ),
    .mOutC_tvalid     (m2C_tvalid   ),
    .mOutC_tdata      (m2C_tdata    ),
    .sInAT_tready     (s2AT_tready  ),
    .sInAT_tvalid     (s2AT_tvalid  ),
    .sInAT_tdata      (s2AT_tdata   ),
    .sInBT_tready     (s2BT_tready  ),
    .sInBT_tvalid     (s2BT_tvalid  ),
    .sInBT_tdata      (s2BT_tdata   ),
    .mOutCT_tready    (m2CT_tready  ),
    .mOutCT_tvalid    (m2CT_tvalid  ),
    .mOutCT_tdata     (m2CT_tdata   ),
    .scInA_tready     (w2cA_tready  ),
    .scInA_tvalid     (w2cA_tvalid  ),
    .scInA_tdata      (w2cA_tdata   ),
    .scInB_tready     (w2cB_tready  ),
    .scInB_tvalid     (w2cB_tvalid  ),
    .scInB_tdata      (w2cB_tdata   ),
    .mcOutC_tready    (w2cC_tready  ),
    .mcOutC_tvalid    (w2cC_tvalid  ),
    .mcOutC_tdata     (w2cC_tdata   ),
    .sAccInC_tready   (s2C_tready   ),
    .sAccInC_tvalid   (s2C_tvalid   ),
    .sAccInC_tdata    (s2C_tdata    ),
    .mAccOutA_tready  (m2A_tready   ),
    .mAccOutA_tvalid  (m2A_tvalid   ),
    .mAccOutA_tdata   (m2A_tdata    ),
    .mAccOutB_tready  (m2B_tready   ),
    .mAccOutB_tvalid  (m2B_tvalid   ),
    .mAccOutB_tdata   (m2B_tdata    ),
    .CONF             (acc2_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc3_couple (
    .sInA_tready      (s3A_tready   ),
    .sInA_tvalid      (s3A_tvalid   ),
    .sInA_tdata       (s3A_tdata    ),
    .sInB_tready      (s3B_tready   ),
    .sInB_tvalid      (s3B_tvalid   ),
    .sInB_tdata       (s3B_tdata    ),
    .mOutC_tready     (m3C_tready   ),
    .mOutC_tvalid     (m3C_tvalid   ),
    .mOutC_tdata      (m3C_tdata    ),
    .sInAT_tready     (s3AT_tready  ),
    .sInAT_tvalid     (s3AT_tvalid  ),
    .sInAT_tdata      (s3AT_tdata   ),
    .sInBT_tready     (s3BT_tready  ),
    .sInBT_tvalid     (s3BT_tvalid  ),
    .sInBT_tdata      (s3BT_tdata   ),
    .mOutCT_tready    (m3CT_tready  ),
    .mOutCT_tvalid    (m3CT_tvalid  ),
    .mOutCT_tdata     (m3CT_tdata   ),
    .scInA_tready     (w3cA_tready  ),
    .scInA_tvalid     (w3cA_tvalid  ),
    .scInA_tdata      (w3cA_tdata   ),
    .scInB_tready     (w3cB_tready  ),
    .scInB_tvalid     (w3cB_tvalid  ),
    .scInB_tdata      (w3cB_tdata   ),
    .mcOutC_tready    (w3cC_tready  ),
    .mcOutC_tvalid    (w3cC_tvalid  ),
    .mcOutC_tdata     (w3cC_tdata   ),
    .sAccInC_tready   (s3C_tready   ),
    .sAccInC_tvalid   (s3C_tvalid   ),
    .sAccInC_tdata    (s3C_tdata    ),
    .mAccOutA_tready  (m3A_tready   ),
    .mAccOutA_tvalid  (m3A_tvalid   ),
    .mAccOutA_tdata   (m3A_tdata    ),
    .mAccOutB_tready  (m3B_tready   ),
    .mAccOutB_tvalid  (m3B_tvalid   ),
    .mAccOutB_tdata   (m3B_tdata    ),
    .CONF             (acc3_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc4_couple (
    .sInA_tready      (s4A_tready   ),
    .sInA_tvalid      (s4A_tvalid   ),
    .sInA_tdata       (s4A_tdata    ),
    .sInB_tready      (s4B_tready   ),
    .sInB_tvalid      (s4B_tvalid   ),
    .sInB_tdata       (s4B_tdata    ),
    .mOutC_tready     (m4C_tready   ),
    .mOutC_tvalid     (m4C_tvalid   ),
    .mOutC_tdata      (m4C_tdata    ),
    .sInAT_tready     (s4AT_tready  ),
    .sInAT_tvalid     (s4AT_tvalid  ),
    .sInAT_tdata      (s4AT_tdata   ),
    .sInBT_tready     (s4BT_tready  ),
    .sInBT_tvalid     (s4BT_tvalid  ),
    .sInBT_tdata      (s4BT_tdata   ),
    .mOutCT_tready    (m4CT_tready  ),
    .mOutCT_tvalid    (m4CT_tvalid  ),
    .mOutCT_tdata     (m4CT_tdata   ),
    .scInA_tready     (w4cA_tready  ),
    .scInA_tvalid     (w4cA_tvalid  ),
    .scInA_tdata      (w4cA_tdata   ),
    .scInB_tready     (w4cB_tready  ),
    .scInB_tvalid     (w4cB_tvalid  ),
    .scInB_tdata      (w4cB_tdata   ),
    .mcOutC_tready    (w4cC_tready  ),
    .mcOutC_tvalid    (w4cC_tvalid  ),
    .mcOutC_tdata     (w4cC_tdata   ),
    .sAccInC_tready   (s4C_tready   ),
    .sAccInC_tvalid   (s4C_tvalid   ),
    .sAccInC_tdata    (s4C_tdata    ),
    .mAccOutA_tready  (m4A_tready   ),
    .mAccOutA_tvalid  (m4A_tvalid   ),
    .mAccOutA_tdata   (m4A_tdata    ),
    .mAccOutB_tready  (m4B_tready   ),
    .mAccOutB_tvalid  (m4B_tvalid   ),
    .mAccOutB_tdata   (m4B_tdata    ),
    .CONF             (acc4_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_crossbar #(NUM_ACCs) u_crossbar (
    .CONF1_A       (acc1_A1         ),
    .CONF1_B       (acc1_B1         ),
    .sC1_tready    (w1cC_tready     ),
    .sC1_tvalid    (w1cC_tvalid     ),
    .sC1_tdata     (w1cC_tdata      ),
    .mA1_tready    (w1cA_tready     ),
    .mA1_tvalid    (w1cA_tvalid     ),
    .mA1_tdata     (w1cA_tdata      ),
    .mB1_tready    (w1cB_tready     ),
    .mB1_tvalid    (w1cB_tvalid     ),
    .mB1_tdata     (w1cB_tdata      ),
    .CONF2_A       (acc2_A1         ),
    .CONF2_B       (acc2_B1         ),
    .sC2_tready    (w2cC_tready     ),
    .sC2_tvalid    (w2cC_tvalid     ),
    .sC2_tdata     (w2cC_tdata      ),
    .mA2_tready    (w2cA_tready     ),
    .mA2_tvalid    (w2cA_tvalid     ),
    .mA2_tdata     (w2cA_tdata      ),
    .mB2_tready    (w2cB_tready     ),
    .mB2_tvalid    (w2cB_tvalid     ),
    .mB2_tdata     (w2cB_tdata      ),
    .CONF3_A       (acc3_A1         ),
    .CONF3_B       (acc3_B1         ),
    .sC3_tready    (w3cC_tready     ),
    .sC3_tvalid    (w3cC_tvalid     ),
    .sC3_tdata     (w3cC_tdata      ),
    .mA3_tready    (w3cA_tready     ),
    .mA3_tvalid    (w3cA_tvalid     ),
    .mA3_tdata     (w3cA_tdata      ),
    .mB3_tready    (w3cB_tready     ),
    .mB3_tvalid    (w3cB_tvalid     ),
    .mB3_tdata     (w3cB_tdata      ),
    .CONF4_A       (acc4_A1         ),
    .CONF4_B       (acc4_B1         ),
    .sC4_tready    (w4cC_tready     ),
    .sC4_tvalid    (w4cC_tvalid     ),
    .sC4_tdata     (w4cC_tdata      ),
    .mA4_tready    (w4cA_tready     ),
    .mA4_tvalid    (w4cA_tvalid     ),
    .mA4_tdata     (w4cA_tdata      ),
    .mB4_tready    (w4cB_tready     ),
    .mB4_tvalid    (w4cB_tvalid     ),
    .mB4_tdata     (w4cB_tdata      ),
    .CONF5_A       (acc5_A1         ),
    .CONF5_B       (acc5_B1         ),
    .sC5_tready    (w5cC_tready     ),
    .sC5_tvalid    ( 1'd0           ),
    .sC5_tdata     (32'd0           ),
    .mA5_tready    ( 1'd0           ),
    .mA5_tvalid    (w5cA_tvalid     ),
    .mA5_tdata     (w5cA_tdata      ),
    .mB5_tready    ( 1'd0           ),
    .mB5_tvalid    (w5cB_tvalid     ),
    .mB5_tdata     (w5cB_tdata      ),
    .CONF6_A       (acc6_A1         ),
    .CONF6_B       (acc6_B1         ),
    .sC6_tready    (w6cC_tready     ),
    .sC6_tvalid    ( 1'd0           ),
    .sC6_tdata     (32'd0           ),
    .mA6_tready    ( 1'd0           ),
    .mA6_tvalid    (w6cA_tvalid     ),
    .mA6_tdata     (w6cA_tdata      ),
    .mB6_tready    ( 1'd0           ),
    .mB6_tvalid    (w6cB_tvalid     ),
    .mB6_tdata     (w6cB_tdata      ),
    .CONF7_A       (acc7_A1         ),
    .CONF7_B       (acc7_B1         ),
    .sC7_tready    (w7cC_tready     ),
    .sC7_tvalid    ( 1'd0           ),
    .sC7_tdata     (32'd0           ),
    .mA7_tready    ( 1'd0           ),
    .mA7_tvalid    (w7cA_tvalid     ),
    .mA7_tdata     (w7cA_tdata      ),
    .mB7_tready    ( 1'd0           ),
    .mB7_tvalid    (w7cB_tvalid     ),
    .mB7_tdata     (w7cB_tdata      ),
    .CONF8_A       (acc8_A1         ),
    .CONF8_B       (acc8_B1         ),
    .sC8_tready    (w8cC_tready     ),
    .sC8_tvalid    ( 1'd0           ),
    .sC8_tdata     (32'd0           ),
    .mA8_tready    ( 1'd0           ),
    .mA8_tvalid    (w8cA_tvalid     ),
    .mA8_tdata     (w8cA_tdata      ),
    .mB8_tready    ( 1'd0           ),
    .mB8_tvalid    (w8cB_tvalid     ),
    .mB8_tdata     (w8cB_tdata      ),
    .ACLK          (ACLK            ),
    .ARESETN       (ARESETN         )
  );

  jit_dispatch #(NUM_ACCs) u_dispatch(
    .sR_tready     (sCMD_tready     ),
    .sR_tvalid     (sCMD_tvalid     ),
    .sR_tdata      (sCMD_tdata      ),
//  .mR_tready     (mRSP_tready     ),
//  .mR_tvalid     (mRSP_tvalid     ),
//  .mR_tdata      (mRSP_tdata      ),
    .acc1_A1       (acc1_A1         ),
    .acc1_B1       (acc1_B1         ),
    .acc1_C1       (acc1_C1         ),
    .acc1_R1       (ap1_arg1_V      ),
    .acc1_R2       (ap1_arg2_V      ),
    .acc1_R3       (ap1_arg3_V      ),
//  .acc1_done     (ap1_done        ),
//  .acc1_idle     (ap1_idle        ),
//  .acc1_ready    (ap1_ready       ),
//  .acc1_start    (ap1_start       ),
    .acc2_A1       (acc2_A1         ),
    .acc2_B1       (acc2_B1         ),
    .acc2_C1       (acc2_C1         ),
    .acc2_R1       (ap2_arg1_V      ),
    .acc2_R2       (ap2_arg2_V      ),
    .acc2_R3       (ap2_arg3_V      ),
//  .acc2_done     (ap2_done        ),
//  .acc2_idle     (ap2_idle        ),
//  .acc2_ready    (ap2_ready       ),
//  .acc2_start    (ap2_start       ),
    .acc3_A1       (acc3_A1         ),
    .acc3_B1       (acc3_B1         ),
    .acc3_C1       (acc3_C1         ),
    .acc3_R1       (ap3_arg1_V      ),
    .acc3_R2       (ap3_arg2_V      ),
    .acc3_R3       (ap3_arg3_V      ),
//  .acc3_done     (ap3_done        ),
//  .acc3_idle     (ap3_idle        ),
//  .acc3_ready    (ap3_ready       ),
//  .acc3_start    (ap3_start       ),
    .acc4_A1       (acc4_A1         ),
    .acc4_B1       (acc4_B1         ),
    .acc4_C1       (acc4_C1         ),
    .acc4_R1       (ap4_arg1_V      ),
    .acc4_R2       (ap4_arg2_V      ),
    .acc4_R3       (ap4_arg3_V      ),
//  .acc4_done     (ap4_done        ),
//  .acc4_idle     (ap4_idle        ),
//  .acc4_ready    (ap4_ready       ),
//  .acc4_start    (ap4_start       ),
    .acc5_A1       (acc5_A1         ),
    .acc5_B1       (acc5_B1         ),
    .acc5_C1       (acc5_C1         ),
    .acc5_R1       (ap5_arg1_V      ),
    .acc5_R2       (ap5_arg2_V      ),
    .acc5_R3       (ap5_arg3_V      ),
//  .acc5_done     (ap5_done        ),
//  .acc5_idle     (ap5_idle        ),
//  .acc5_ready    (ap5_ready       ),
//  .acc5_start    (ap5_start       ),
    .acc6_A1       (acc6_A1         ),
    .acc6_B1       (acc6_B1         ),
    .acc6_C1       (acc6_C1         ),
    .acc6_R1       (ap6_arg1_V      ),
    .acc6_R2       (ap6_arg2_V      ),
    .acc6_R3       (ap6_arg3_V      ),
//  .acc6_done     (ap6_done        ),
//  .acc6_idle     (ap6_idle        ),
//  .acc6_ready    (ap6_ready       ),
//  .acc6_start    (ap6_start       ),
    .acc7_A1       (acc7_A1         ),
    .acc7_B1       (acc7_B1         ),
    .acc7_C1       (acc7_C1         ),
    .acc7_R1       (ap7_arg1_V      ),
    .acc7_R2       (ap7_arg2_V      ),
    .acc7_R3       (ap7_arg3_V      ),
//  .acc7_done     (ap7_done        ),
//  .acc7_idle     (ap7_idle        ),
//  .acc7_ready    (ap7_ready       ),
//  .acc7_start    (ap7_start       ),
    .acc8_A1       (acc8_A1         ),
    .acc8_B1       (acc8_B1         ),
    .acc8_C1       (acc8_C1         ),
    .acc8_R1       (ap8_arg1_V      ),
    .acc8_R2       (ap8_arg2_V      ),
    .acc8_R3       (ap8_arg3_V      ),
//  .acc8_done     (ap8_done        ),
//  .acc8_idle     (ap8_idle        ),
//  .acc8_ready    (ap8_ready       ),
//  .acc8_start    (ap8_start       ),
    .ACLK          (ACLK            ),
    .ARESETN       (ARESETN         )
  );

end
endgenerate // NUM_ACCs == 8
//       _    ____ ____            ___
//      / \  / ___/ ___|___   _   ( _ )
//     / _ \| |  | |   / __| (_)  / _ \
//    / ___ \ |__| |___\__ \  _  | (_) |
//   /_/   \_\____\____|___/ (_)  \___/
//
generate if (NUM_ACCs == 8) begin

  jit_couple u_acc1_couple (
    .sInA_tready      (s1A_tready   ),
    .sInA_tvalid      (s1A_tvalid   ),
    .sInA_tdata       (s1A_tdata    ),
    .sInB_tready      (s1B_tready   ),
    .sInB_tvalid      (s1B_tvalid   ),
    .sInB_tdata       (s1B_tdata    ),
    .mOutC_tready     (m1C_tready   ),
    .mOutC_tvalid     (m1C_tvalid   ),
    .mOutC_tdata      (m1C_tdata    ),
    .sInAT_tready     (s1AT_tready  ),
    .sInAT_tvalid     (s1AT_tvalid  ),
    .sInAT_tdata      (s1AT_tdata   ),
    .sInBT_tready     (s1BT_tready  ),
    .sInBT_tvalid     (s1BT_tvalid  ),
    .sInBT_tdata      (s1BT_tdata   ),
    .mOutCT_tready    (m1CT_tready  ),
    .mOutCT_tvalid    (m1CT_tvalid  ),
    .mOutCT_tdata     (m1CT_tdata   ),
    .scInA_tready     (w1cA_tready  ),
    .scInA_tvalid     (w1cA_tvalid  ),
    .scInA_tdata      (w1cA_tdata   ),
    .scInB_tready     (w1cB_tready  ),
    .scInB_tvalid     (w1cB_tvalid  ),
    .scInB_tdata      (w1cB_tdata   ),
    .mcOutC_tready    (w1cC_tready  ),
    .mcOutC_tvalid    (w1cC_tvalid  ),
    .mcOutC_tdata     (w1cC_tdata   ),
    .sAccInC_tready   (s1C_tready   ),
    .sAccInC_tvalid   (s1C_tvalid   ),
    .sAccInC_tdata    (s1C_tdata    ),
    .mAccOutA_tready  (m1A_tready   ),
    .mAccOutA_tvalid  (m1A_tvalid   ),
    .mAccOutA_tdata   (m1A_tdata    ),
    .mAccOutB_tready  (m1B_tready   ),
    .mAccOutB_tvalid  (m1B_tvalid   ),
    .mAccOutB_tdata   (m1B_tdata    ),
    .CONF             (acc1_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc2_couple (
    .sInA_tready      (s2A_tready   ),
    .sInA_tvalid      (s2A_tvalid   ),
    .sInA_tdata       (s2A_tdata    ),
    .sInB_tready      (s2B_tready   ),
    .sInB_tvalid      (s2B_tvalid   ),
    .sInB_tdata       (s2B_tdata    ),
    .mOutC_tready     (m2C_tready   ),
    .mOutC_tvalid     (m2C_tvalid   ),
    .mOutC_tdata      (m2C_tdata    ),
    .sInAT_tready     (s2AT_tready  ),
    .sInAT_tvalid     (s2AT_tvalid  ),
    .sInAT_tdata      (s2AT_tdata   ),
    .sInBT_tready     (s2BT_tready  ),
    .sInBT_tvalid     (s2BT_tvalid  ),
    .sInBT_tdata      (s2BT_tdata   ),
    .mOutCT_tready    (m2CT_tready  ),
    .mOutCT_tvalid    (m2CT_tvalid  ),
    .mOutCT_tdata     (m2CT_tdata   ),
    .scInA_tready     (w2cA_tready  ),
    .scInA_tvalid     (w2cA_tvalid  ),
    .scInA_tdata      (w2cA_tdata   ),
    .scInB_tready     (w2cB_tready  ),
    .scInB_tvalid     (w2cB_tvalid  ),
    .scInB_tdata      (w2cB_tdata   ),
    .mcOutC_tready    (w2cC_tready  ),
    .mcOutC_tvalid    (w2cC_tvalid  ),
    .mcOutC_tdata     (w2cC_tdata   ),
    .sAccInC_tready   (s2C_tready   ),
    .sAccInC_tvalid   (s2C_tvalid   ),
    .sAccInC_tdata    (s2C_tdata    ),
    .mAccOutA_tready  (m2A_tready   ),
    .mAccOutA_tvalid  (m2A_tvalid   ),
    .mAccOutA_tdata   (m2A_tdata    ),
    .mAccOutB_tready  (m2B_tready   ),
    .mAccOutB_tvalid  (m2B_tvalid   ),
    .mAccOutB_tdata   (m2B_tdata    ),
    .CONF             (acc2_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc3_couple (
    .sInA_tready      (s3A_tready   ),
    .sInA_tvalid      (s3A_tvalid   ),
    .sInA_tdata       (s3A_tdata    ),
    .sInB_tready      (s3B_tready   ),
    .sInB_tvalid      (s3B_tvalid   ),
    .sInB_tdata       (s3B_tdata    ),
    .mOutC_tready     (m3C_tready   ),
    .mOutC_tvalid     (m3C_tvalid   ),
    .mOutC_tdata      (m3C_tdata    ),
    .sInAT_tready     (s3AT_tready  ),
    .sInAT_tvalid     (s3AT_tvalid  ),
    .sInAT_tdata      (s3AT_tdata   ),
    .sInBT_tready     (s3BT_tready  ),
    .sInBT_tvalid     (s3BT_tvalid  ),
    .sInBT_tdata      (s3BT_tdata   ),
    .mOutCT_tready    (m3CT_tready  ),
    .mOutCT_tvalid    (m3CT_tvalid  ),
    .mOutCT_tdata     (m3CT_tdata   ),
    .scInA_tready     (w3cA_tready  ),
    .scInA_tvalid     (w3cA_tvalid  ),
    .scInA_tdata      (w3cA_tdata   ),
    .scInB_tready     (w3cB_tready  ),
    .scInB_tvalid     (w3cB_tvalid  ),
    .scInB_tdata      (w3cB_tdata   ),
    .mcOutC_tready    (w3cC_tready  ),
    .mcOutC_tvalid    (w3cC_tvalid  ),
    .mcOutC_tdata     (w3cC_tdata   ),
    .sAccInC_tready   (s3C_tready   ),
    .sAccInC_tvalid   (s3C_tvalid   ),
    .sAccInC_tdata    (s3C_tdata    ),
    .mAccOutA_tready  (m3A_tready   ),
    .mAccOutA_tvalid  (m3A_tvalid   ),
    .mAccOutA_tdata   (m3A_tdata    ),
    .mAccOutB_tready  (m3B_tready   ),
    .mAccOutB_tvalid  (m3B_tvalid   ),
    .mAccOutB_tdata   (m3B_tdata    ),
    .CONF             (acc3_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc4_couple (
    .sInA_tready      (s4A_tready   ),
    .sInA_tvalid      (s4A_tvalid   ),
    .sInA_tdata       (s4A_tdata    ),
    .sInB_tready      (s4B_tready   ),
    .sInB_tvalid      (s4B_tvalid   ),
    .sInB_tdata       (s4B_tdata    ),
    .mOutC_tready     (m4C_tready   ),
    .mOutC_tvalid     (m4C_tvalid   ),
    .mOutC_tdata      (m4C_tdata    ),
    .sInAT_tready     (s4AT_tready  ),
    .sInAT_tvalid     (s4AT_tvalid  ),
    .sInAT_tdata      (s4AT_tdata   ),
    .sInBT_tready     (s4BT_tready  ),
    .sInBT_tvalid     (s4BT_tvalid  ),
    .sInBT_tdata      (s4BT_tdata   ),
    .mOutCT_tready    (m4CT_tready  ),
    .mOutCT_tvalid    (m4CT_tvalid  ),
    .mOutCT_tdata     (m4CT_tdata   ),
    .scInA_tready     (w4cA_tready  ),
    .scInA_tvalid     (w4cA_tvalid  ),
    .scInA_tdata      (w4cA_tdata   ),
    .scInB_tready     (w4cB_tready  ),
    .scInB_tvalid     (w4cB_tvalid  ),
    .scInB_tdata      (w4cB_tdata   ),
    .mcOutC_tready    (w4cC_tready  ),
    .mcOutC_tvalid    (w4cC_tvalid  ),
    .mcOutC_tdata     (w4cC_tdata   ),
    .sAccInC_tready   (s4C_tready   ),
    .sAccInC_tvalid   (s4C_tvalid   ),
    .sAccInC_tdata    (s4C_tdata    ),
    .mAccOutA_tready  (m4A_tready   ),
    .mAccOutA_tvalid  (m4A_tvalid   ),
    .mAccOutA_tdata   (m4A_tdata    ),
    .mAccOutB_tready  (m4B_tready   ),
    .mAccOutB_tvalid  (m4B_tvalid   ),
    .mAccOutB_tdata   (m4B_tdata    ),
    .CONF             (acc4_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc5_couple (
    .sInA_tready      (s5A_tready   ),
    .sInA_tvalid      (s5A_tvalid   ),
    .sInA_tdata       (s5A_tdata    ),
    .sInB_tready      (s5B_tready   ),
    .sInB_tvalid      (s5B_tvalid   ),
    .sInB_tdata       (s5B_tdata    ),
    .mOutC_tready     (m5C_tready   ),
    .mOutC_tvalid     (m5C_tvalid   ),
    .mOutC_tdata      (m5C_tdata    ),
    .sInAT_tready     (s5AT_tready  ),
    .sInAT_tvalid     (s5AT_tvalid  ),
    .sInAT_tdata      (s5AT_tdata   ),
    .sInBT_tready     (s5BT_tready  ),
    .sInBT_tvalid     (s5BT_tvalid  ),
    .sInBT_tdata      (s5BT_tdata   ),
    .mOutCT_tready    (m5CT_tready  ),
    .mOutCT_tvalid    (m5CT_tvalid  ),
    .mOutCT_tdata     (m5CT_tdata   ),
    .scInA_tready     (w5cA_tready  ),
    .scInA_tvalid     (w5cA_tvalid  ),
    .scInA_tdata      (w5cA_tdata   ),
    .scInB_tready     (w5cB_tready  ),
    .scInB_tvalid     (w5cB_tvalid  ),
    .scInB_tdata      (w5cB_tdata   ),
    .mcOutC_tready    (w5cC_tready  ),
    .mcOutC_tvalid    (w5cC_tvalid  ),
    .mcOutC_tdata     (w5cC_tdata   ),
    .sAccInC_tready   (s5C_tready   ),
    .sAccInC_tvalid   (s5C_tvalid   ),
    .sAccInC_tdata    (s5C_tdata    ),
    .mAccOutA_tready  (m5A_tready   ),
    .mAccOutA_tvalid  (m5A_tvalid   ),
    .mAccOutA_tdata   (m5A_tdata    ),
    .mAccOutB_tready  (m5B_tready   ),
    .mAccOutB_tvalid  (m5B_tvalid   ),
    .mAccOutB_tdata   (m5B_tdata    ),
    .CONF             (acc5_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple       u_acc6_couple (
    .sInA_tready      (s6A_tready   ),
    .sInA_tvalid      (s6A_tvalid   ),
    .sInA_tdata       (s6A_tdata    ),
    .sInB_tready      (s6B_tready   ),
    .sInB_tvalid      (s6B_tvalid   ),
    .sInB_tdata       (s6B_tdata    ),
    .mOutC_tready     (m6C_tready   ),
    .mOutC_tvalid     (m6C_tvalid   ),
    .mOutC_tdata      (m6C_tdata    ),
    .sInAT_tready     (s6AT_tready  ),
    .sInAT_tvalid     (s6AT_tvalid  ),
    .sInAT_tdata      (s6AT_tdata   ),
    .sInBT_tready     (s6BT_tready  ),
    .sInBT_tvalid     (s6BT_tvalid  ),
    .sInBT_tdata      (s6BT_tdata   ),
    .mOutCT_tready    (m6CT_tready  ),
    .mOutCT_tvalid    (m6CT_tvalid  ),
    .mOutCT_tdata     (m6CT_tdata   ),
    .scInA_tready     (w6cA_tready  ),
    .scInA_tvalid     (w6cA_tvalid  ),
    .scInA_tdata      (w6cA_tdata   ),
    .scInB_tready     (w6cB_tready  ),
    .scInB_tvalid     (w6cB_tvalid  ),
    .scInB_tdata      (w6cB_tdata   ),
    .mcOutC_tready    (w6cC_tready  ),
    .mcOutC_tvalid    (w6cC_tvalid  ),
    .mcOutC_tdata     (w6cC_tdata   ),
    .sAccInC_tready   (s6C_tready   ),
    .sAccInC_tvalid   (s6C_tvalid   ),
    .sAccInC_tdata    (s6C_tdata    ),
    .mAccOutA_tready  (m6A_tready   ),
    .mAccOutA_tvalid  (m6A_tvalid   ),
    .mAccOutA_tdata   (m6A_tdata    ),
    .mAccOutB_tready  (m6B_tready   ),
    .mAccOutB_tvalid  (m6B_tvalid   ),
    .mAccOutB_tdata   (m6B_tdata    ),
    .CONF             (acc6_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc7_couple (
    .sInA_tready      (s7A_tready   ),
    .sInA_tvalid      (s7A_tvalid   ),
    .sInA_tdata       (s7A_tdata    ),
    .sInB_tready      (s7B_tready   ),
    .sInB_tvalid      (s7B_tvalid   ),
    .sInB_tdata       (s7B_tdata    ),
    .mOutC_tready     (m7C_tready   ),
    .mOutC_tvalid     (m7C_tvalid   ),
    .mOutC_tdata      (m7C_tdata    ),
    .sInAT_tready     (s7AT_tready  ),
    .sInAT_tvalid     (s7AT_tvalid  ),
    .sInAT_tdata      (s7AT_tdata   ),
    .sInBT_tready     (s7BT_tready  ),
    .sInBT_tvalid     (s7BT_tvalid  ),
    .sInBT_tdata      (s7BT_tdata   ),
    .mOutCT_tready    (m7CT_tready  ),
    .mOutCT_tvalid    (m7CT_tvalid  ),
    .mOutCT_tdata     (m7CT_tdata   ),
    .scInA_tready     (w7cA_tready  ),
    .scInA_tvalid     (w7cA_tvalid  ),
    .scInA_tdata      (w7cA_tdata   ),
    .scInB_tready     (w7cB_tready  ),
    .scInB_tvalid     (w7cB_tvalid  ),
    .scInB_tdata      (w7cB_tdata   ),
    .mcOutC_tready    (w7cC_tready  ),
    .mcOutC_tvalid    (w7cC_tvalid  ),
    .mcOutC_tdata     (w7cC_tdata   ),
    .sAccInC_tready   (s7C_tready   ),
    .sAccInC_tvalid   (s7C_tvalid   ),
    .sAccInC_tdata    (s7C_tdata    ),
    .mAccOutA_tready  (m7A_tready   ),
    .mAccOutA_tvalid  (m7A_tvalid   ),
    .mAccOutA_tdata   (m7A_tdata    ),
    .mAccOutB_tready  (m7B_tready   ),
    .mAccOutB_tvalid  (m7B_tvalid   ),
    .mAccOutB_tdata   (m7B_tdata    ),
    .CONF             (acc7_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_couple u_acc8_couple (
    .sInA_tready      (s8A_tready   ),
    .sInA_tvalid      (s8A_tvalid   ),
    .sInA_tdata       (s8A_tdata    ),
    .sInB_tready      (s8B_tready   ),
    .sInB_tvalid      (s8B_tvalid   ),
    .sInB_tdata       (s8B_tdata    ),
    .mOutC_tready     (m8C_tready   ),
    .mOutC_tvalid     (m8C_tvalid   ),
    .mOutC_tdata      (m8C_tdata    ),
    .sInAT_tready     (s8AT_tready  ),
    .sInAT_tvalid     (s8AT_tvalid  ),
    .sInAT_tdata      (s8AT_tdata   ),
    .sInBT_tready     (s8BT_tready  ),
    .sInBT_tvalid     (s8BT_tvalid  ),
    .sInBT_tdata      (s8BT_tdata   ),
    .mOutCT_tready    (m8CT_tready  ),
    .mOutCT_tvalid    (m8CT_tvalid  ),
    .mOutCT_tdata     (m8CT_tdata   ),
    .scInA_tready     (w8cA_tready  ),
    .scInA_tvalid     (w8cA_tvalid  ),
    .scInA_tdata      (w8cA_tdata   ),
    .scInB_tready     (w8cB_tready  ),
    .scInB_tvalid     (w8cB_tvalid  ),
    .scInB_tdata      (w8cB_tdata   ),
    .mcOutC_tready    (w8cC_tready  ),
    .mcOutC_tvalid    (w8cC_tvalid  ),
    .mcOutC_tdata     (w8cC_tdata   ),
    .sAccInC_tready   (s8C_tready   ),
    .sAccInC_tvalid   (s8C_tvalid   ),
    .sAccInC_tdata    (s8C_tdata    ),
    .mAccOutA_tready  (m8A_tready   ),
    .mAccOutA_tvalid  (m8A_tvalid   ),
    .mAccOutA_tdata   (m8A_tdata    ),
    .mAccOutB_tready  (m8B_tready   ),
    .mAccOutB_tvalid  (m8B_tvalid   ),
    .mAccOutB_tdata   (m8B_tdata    ),
    .CONF             (acc8_C1      ),
    .ACLK             (ACLK         ),
    .ARESETN          (ARESETN      )
  );

  jit_crossbar #(NUM_ACCs) u_crossbar (
    .CONF1_A       (acc1_A1         ),
    .CONF1_B       (acc1_B1         ),
    .sC1_tready    (w1cC_tready     ),
    .sC1_tvalid    (w1cC_tvalid     ),
    .sC1_tdata     (w1cC_tdata      ),
    .mA1_tready    (w1cA_tready     ),
    .mA1_tvalid    (w1cA_tvalid     ),
    .mA1_tdata     (w1cA_tdata      ),
    .mB1_tready    (w1cB_tready     ),
    .mB1_tvalid    (w1cB_tvalid     ),
    .mB1_tdata     (w1cB_tdata      ),
    .CONF2_A       (acc2_A1         ),
    .CONF2_B       (acc2_B1         ),
    .sC2_tready    (w2cC_tready     ),
    .sC2_tvalid    (w2cC_tvalid     ),
    .sC2_tdata     (w2cC_tdata      ),
    .mA2_tready    (w2cA_tready     ),
    .mA2_tvalid    (w2cA_tvalid     ),
    .mA2_tdata     (w2cA_tdata      ),
    .mB2_tready    (w2cB_tready     ),
    .mB2_tvalid    (w2cB_tvalid     ),
    .mB2_tdata     (w2cB_tdata      ),
    .CONF3_A       (acc3_A1         ),
    .CONF3_B       (acc3_B1         ),
    .sC3_tready    (w3cC_tready     ),
    .sC3_tvalid    (w3cC_tvalid     ),
    .sC3_tdata     (w3cC_tdata      ),
    .mA3_tready    (w3cA_tready     ),
    .mA3_tvalid    (w3cA_tvalid     ),
    .mA3_tdata     (w3cA_tdata      ),
    .mB3_tready    (w3cB_tready     ),
    .mB3_tvalid    (w3cB_tvalid     ),
    .mB3_tdata     (w3cB_tdata      ),
    .CONF4_A       (acc4_A1         ),
    .CONF4_B       (acc4_B1         ),
    .sC4_tready    (w4cC_tready     ),
    .sC4_tvalid    (w4cC_tvalid     ),
    .sC4_tdata     (w4cC_tdata      ),
    .mA4_tready    (w4cA_tready     ),
    .mA4_tvalid    (w4cA_tvalid     ),
    .mA4_tdata     (w4cA_tdata      ),
    .mB4_tready    (w4cB_tready     ),
    .mB4_tvalid    (w4cB_tvalid     ),
    .mB4_tdata     (w4cB_tdata      ),
    .CONF5_A       (acc5_A1         ),
    .CONF5_B       (acc5_B1         ),
    .sC5_tready    (w5cC_tready     ),
    .sC5_tvalid    (w5cC_tvalid     ),
    .sC5_tdata     (w5cC_tdata      ),
    .mA5_tready    (w5cA_tready     ),
    .mA5_tvalid    (w5cA_tvalid     ),
    .mA5_tdata     (w5cA_tdata      ),
    .mB5_tready    (w5cB_tready     ),
    .mB5_tvalid    (w5cB_tvalid     ),
    .mB5_tdata     (w5cB_tdata      ),
    .CONF6_A       (acc6_A1         ),
    .CONF6_B       (acc6_B1         ),
    .sC6_tready    (w6cC_tready     ),
    .sC6_tvalid    (w6cC_tvalid     ),
    .sC6_tdata     (w6cC_tdata      ),
    .mA6_tready    (w6cA_tready     ),
    .mA6_tvalid    (w6cA_tvalid     ),
    .mA6_tdata     (w6cA_tdata      ),
    .mB6_tready    (w6cB_tready     ),
    .mB6_tvalid    (w6cB_tvalid     ),
    .mB6_tdata     (w6cB_tdata      ),
    .CONF7_A       (acc7_A1         ),
    .CONF7_B       (acc7_B1         ),
    .sC7_tready    (w7cC_tready     ),
    .sC7_tvalid    (w7cC_tvalid     ),
    .sC7_tdata     (w7cC_tdata      ),
    .mA7_tready    (w7cA_tready     ),
    .mA7_tvalid    (w7cA_tvalid     ),
    .mA7_tdata     (w7cA_tdata      ),
    .mB7_tready    (w7cB_tready     ),
    .mB7_tvalid    (w7cB_tvalid     ),
    .mB7_tdata     (w7cB_tdata      ),
    .CONF8_A       (acc8_A1         ),
    .CONF8_B       (acc8_B1         ),
    .sC8_tready    (w8cC_tready     ),
    .sC8_tvalid    (w8cC_tvalid     ),
    .sC8_tdata     (w8cC_tdata      ),
    .mA8_tready    (w8cA_tready     ),
    .mA8_tvalid    (w8cA_tvalid     ),
    .mA8_tdata     (w8cA_tdata      ),
    .mB8_tready    (w8cB_tready     ),
    .mB8_tvalid    (w8cB_tvalid     ),
    .mB8_tdata     (w8cB_tdata      ),
    .ACLK          (ACLK            ),
    .ARESETN       (ARESETN         )
  );

  jit_dispatch #(NUM_ACCs) u_dispatch(
    .sR_tready     (sCMD_tready     ),
    .sR_tvalid     (sCMD_tvalid     ),
    .sR_tdata      (sCMD_tdata      ),
//  .mR_tready     (mRSP_tready     ),
//  .mR_tvalid     (mRSP_tvalid     ),
//  .mR_tdata      (mRSP_tdata      ),
    .acc1_A1       (acc1_A1         ),
    .acc1_B1       (acc1_B1         ),
    .acc1_C1       (acc1_C1         ),
    .acc1_R1       (ap1_arg1_V      ),
    .acc1_R2       (ap1_arg2_V      ),
    .acc1_R3       (ap1_arg3_V      ),
//  .acc1_done     (ap1_done        ),
//  .acc1_idle     (ap1_idle        ),
//  .acc1_ready    (ap1_ready       ),
//  .acc1_start    (ap1_start       ),
    .acc2_A1       (acc2_A1         ),
    .acc2_B1       (acc2_B1         ),
    .acc2_C1       (acc2_C1         ),
    .acc2_R1       (ap2_arg1_V      ),
    .acc2_R2       (ap2_arg2_V      ),
    .acc2_R3       (ap2_arg3_V      ),
//  .acc2_done     (ap2_done        ),
//  .acc2_idle     (ap2_idle        ),
//  .acc2_ready    (ap2_ready       ),
//  .acc2_start    (ap2_start       ),
    .acc3_A1       (acc3_A1         ),
    .acc3_B1       (acc3_B1         ),
    .acc3_C1       (acc3_C1         ),
    .acc3_R1       (ap3_arg1_V      ),
    .acc3_R2       (ap3_arg2_V      ),
    .acc3_R3       (ap3_arg3_V      ),
//  .acc3_done     (ap3_done        ),
//  .acc3_idle     (ap3_idle        ),
//  .acc3_ready    (ap3_ready       ),
//  .acc3_start    (ap3_start       ),
    .acc4_A1       (acc4_A1         ),
    .acc4_B1       (acc4_B1         ),
    .acc4_C1       (acc4_C1         ),
    .acc4_R1       (ap4_arg1_V      ),
    .acc4_R2       (ap4_arg2_V      ),
    .acc4_R3       (ap4_arg3_V      ),
//  .acc4_done     (ap4_done        ),
//  .acc4_idle     (ap4_idle        ),
//  .acc4_ready    (ap4_ready       ),
//  .acc4_start    (ap4_start       ),
    .acc5_A1       (acc5_A1         ),
    .acc5_B1       (acc5_B1         ),
    .acc5_C1       (acc5_C1         ),
    .acc5_R1       (ap5_arg1_V      ),
    .acc5_R2       (ap5_arg2_V      ),
    .acc5_R3       (ap5_arg3_V      ),
//  .acc5_done     (ap5_done        ),
//  .acc5_idle     (ap5_idle        ),
//  .acc5_ready    (ap5_ready       ),
//  .acc5_start    (ap5_start       ),
    .acc6_A1       (acc6_A1         ),
    .acc6_B1       (acc6_B1         ),
    .acc6_C1       (acc6_C1         ),
    .acc6_R1       (ap6_arg1_V      ),
    .acc6_R2       (ap6_arg2_V      ),
    .acc6_R3       (ap6_arg3_V      ),
//  .acc6_done     (ap6_done        ),
//  .acc6_idle     (ap6_idle        ),
//  .acc6_ready    (ap6_ready       ),
//  .acc6_start    (ap6_start       ),
    .acc7_A1       (acc7_A1         ),
    .acc7_B1       (acc7_B1         ),
    .acc7_C1       (acc7_C1         ),
    .acc7_R1       (ap7_arg1_V      ),
    .acc7_R2       (ap7_arg2_V      ),
    .acc7_R3       (ap7_arg3_V      ),
//  .acc7_done     (ap7_done        ),
//  .acc7_idle     (ap7_idle        ),
//  .acc7_ready    (ap7_ready       ),
//  .acc7_start    (ap7_start       ),
    .acc8_A1       (acc8_A1         ),
    .acc8_B1       (acc8_B1         ),
    .acc8_C1       (acc8_C1         ),
    .acc8_R1       (ap8_arg1_V      ),
    .acc8_R2       (ap8_arg2_V      ),
    .acc8_R3       (ap8_arg3_V      ),
//  .acc8_done     (ap8_done        ),
//  .acc8_idle     (ap8_idle        ),
//  .acc8_ready    (ap8_ready       ),
//  .acc8_start    (ap8_start       ),
    .ACLK          (ACLK            ),
    .ARESETN       (ARESETN         )
  );

end
endgenerate // NUM_ACCs == 8

endmodule
